---  В этом файле приводится описание центрального устройства управления ЦУУ.
-- Оно должно формировать управляющие сигналы для ОП, РП и спроектированного ранее арифметического устройства
-- Внешними сигналами для ЦУУ являются сигналы set, по которому ЦУУ, устанавливается в исходное состояние и тактовый сигнал clk
-- Для арифметического устройства оно готовит операнды А и В, задает сор и подает сигнал начала операции sno, после их подготовки
-- Из арифметического устройства оно забирает результат,
-- для умножения это 2n-разрядное произведение, для сложения -n-разрядная сумма и двухразрядный признак результата.
-- Сигналом, подтверждающим выполнение операции в арифметическом устройстве, является сигнал конца операции sko
-- Для оперативной памяти оно формирует следующие сигналы:
-- data_in_OP [7:0] - данные для записи в ОП
-- address_OP [7:0] - адрес, для обращения к ОП
-- wr_en_OP - сигнал записи в ОП, если этот сигнал не активен ОП выполняет чтение
-- Из ОП в ЦУУ поступает сигнал 
-- data_out_OP [7:0] - данные, считанные из ОП
-- Для регистровой памяти РП ЦУУ формирует следующие сигналы 
-- data_a_RP - данные для записи в РП, через порт а
-- address_a_RP [2:0] - адрес, для обращения к RП, через порт a
-- wren_a_RP - сигнал записи через порт а в РП, если этот сигнал не активен PП выполняет чтение
-- data_b_RP - данные для записи в РП, через порт b
-- address_b_RP [2:0] - адрес, для обращения к RП, через порт b
-- wr_en_b_RP - сигнал записи через порт b в РП, если этот сигнал не активен PП выполняет чтение
-- q_a - данные, считываемые из РП, через порт а
-- q_b - данные, считываемые из РП, через порт b



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.numeric_std.all; -- добавляем библиотеку
LIBRARY work;

--LIBRARY altera_mf;

--USE altera_mf.altera_mf_components.all;

entity Module_CYY is
generic (n:integer:=8);     -- n параметр, задает разрядность операндов
	port
	(	
		clk		 : in	std_logic; -- тактовый сигнал
		set 	 : in	std_logic; --  сигнал начальной установки
		f_com    : buffer std_logic_vector(1 downto 0); -- теперь определяется по команде в RK - УП; 1 - РР; 0 - ПР
-- Для взаимодействия с АУ
		a 			 : out STD_LOGIC_VECTOR (n-1 downto 0);-- первый операнд для АУ		
		b 			 : out STD_LOGIC_VECTOR (n-1 downto 0);-- второй операнд для АУ		
		cop		     : out std_logic; --  код операции 1-умножение,0 - сложение для АУ
		sno		     : out std_logic; -- сигнал начала операции для АУ
		rr 		     : in STD_LOGIC_VECTOR (2*n-1 downto 0);-- результат из АУ
        priznak      : in STD_LOGIC_VECTOR (1 downto 0); -- признак результата из АУ
		sko	 	     : in std_logic; -- сигнал конца операции из АУ
-- Для наблюдения внутренних сигналов во время отладки проекта
		signal RA    : buffer STD_LOGIC_VECTOR (7 downto 0);-- регистр адреса, для адресации операнда в ОП
		signal CK    : buffer STD_LOGIC_VECTOR (7 downto 0);-- счетчик команд, для адресации текущей команды в ОП
		signal RK    : buffer STD_LOGIC_VECTOR (7 downto 0);-- регистр команд, для хранения текущей выполняемой команды
		s_out	     : out STD_LOGIC_VECTOR(2 downto 0);    -- отладочный выход для наблюдения состояний БМК
-- Для взаимодействия с ОП		
		data_in_OP   : out STD_LOGIC_VECTOR (7 downto 0); -- данные для записи в ОП
		address_OP   : out STD_LOGIC_VECTOR (7 downto 0); -- адрес, для обращения к ОП
		wr_en_OP     : out std_logic; -- сигнал записи в ОП, если этот сигнал не активен, ОП выполняет чтение
		data_out_OP  : in  STD_LOGIC_VECTOR (7 downto 0); -- данные, считанные из ОП

-- Для взаимодействия с РП
 		data_a_RP    : out STD_LOGIC_VECTOR (7 downto 0); -- данные для записи в РП, через порт а
		address_a_RP : out STD_LOGIC_VECTOR (2 downto 0); -- адрес, для обращения к RП, через порт a
		wr_en_a_RP 	 : out std_logic; 						  -- сигнал записи через порт а в РП, если этот сигнал не активен PП выполняет чтение
 		data_b_RP 	 : out STD_LOGIC_VECTOR (7 downto 0); -- данные для записи в РП, через порт b
		address_b_RP : out STD_LOGIC_VECTOR (2 downto 0); -- адрес, для обращения к RП, через порт b
  		wr_en_b_RP 	 : out std_logic;					  -- сигнал записи через порт b в РП, если этот сигнал не активен PП выполняет чтение
		q_a 		 : in  STD_LOGIC_VECTOR (7 downto 0);-- данные из РП с порта а	
		q_b 		 : in  STD_LOGIC_VECTOR (7 downto 0) -- данные из РП с порта b
	);

end entity Module_CYY;

architecture arch of Module_CYY is

------------------------------------------------------------------------------------------------------------------------------------------------
-- Декларация сигналов, используемых в проекте 
type state_type is (s0, s1, s2, s3, s4, s5, s6); -- определяем состояния БМК
	signal next_state, state : state_type; -- следующее состояние, текущее состояние
    signal incr_CK	: STD_LOGIC:='0';-- разрешение инкремента СК
    signal summ_CK	: STD_LOGIC:='0';-- вычисление адреса перехода
    signal load_RK	: STD_LOGIC:='0';-- загрузка команды
    signal load_RA	: STD_LOGIC:='0';-- загрузка адреса
    signal IA		: STD_LOGIC_VECTOR (7 downto 0);-- исполнительный адрес операнда в ОП 
    signal incr_RA	: STD_LOGIC:='0';-- разрешение инкремента РА
-----------------------------------------------------------------------------------

begin

-------------------------------------------------------------------------------------------
pr_CK:   process (set, clk) -- этот процесс определяет поведение счетчика команд СК
	
	begin
		if (set='1') then CK<=(others=>'0'); --устанавливаем в начальное состояние
		elsif clk'event and clk='1' then 
		  if (incr_CK='1') then CK<=CK+"00000001"; -- инкремент счетчика
			elsif (summ_CK='1') then CK<= CK+(RK(5)&RK(5)&RK(5 downto 0)); -- вычисление адреса перехода
		  end if;
		 end if;
	end process pr_CK;
---------------------------------------------------------------------------------------	 
pr_RK: process (clk) -- этот процесс определяет поведение регистра команд
	begin
		if clk'event and clk='1' then -- по положительному фронту clk
			if load_RK='1' then -- если есть разрешение на прием команды
			RK<=data_out_OP; -- выполняется прием команды с выхода ОП
			end if;
		end if;
	end process pr_RK;
---------------------------------------------------------------------------------------------
pr_RA: process (clk)-- этот процесс описывает логику работы регистра адреса RA
	begin
		if clk'event and clk='1' then -- по положительному фронту 
		 if load_RA='1' then  RA<=IA; -- если есть разрешение, то загружаем исполнительный адрес первого операнда		
				elsif incr_RA='1' then RA<=RA+1; --инкремент адреса"00000001"
		 end if;
		end if;
end process pr_RA;
------------------------------------------------------------------------------------------------
-- Ниже приводится описание устройства управления для ЦУУ.Реализованы три формата команд ПР,РР и УП
TS: process (clk,set) -- этот процесс определяет текущее состояние МУУ
	 begin
		if set = '1' then
			state <= s0;
		elsif (rising_edge(clk)) then -- по положительному фронту переключаются состояния
			state <= next_state;			
		end if;
	 end process TS;
	 
NS: process (state,set,f_com,sko,priznak) -- этот процесс определяет следующее состояние МУУ, управляющие сигналы
	 begin
-- 

			case state is
				when s0=> -- переходы из s0
				 
					if (set = '0') then
						next_state <= s1; -- если сигнал set не активен,load_RK, incr_CK 
					else
						next_state <= s0; -- иначе состояние не меняется
					end if;
				when s1=>
				   if (f_com = "00") then -- если формат П-Р, то
						next_state <= s2; -- переходим в s2 в случае ПР
					elsif (f_com="01") then
						next_state <= s3; -- переходим в s3 в случае РР
					elsif priznak="10" then
						next_state<=s6;	-- переходим в s6 в случае УП и условие пер выполнено
					else
						next_state<=s0;	-- иначе в s0
					end if;	
				when s2=>
					
						next_state <= s3; -- из s2 всегда переходим в s3 load_RA,

				when s3 =>
						next_state <= s4; -- из s3 всегда переходим в s4, sno=1,summ_RA
						
				when s4 =>
							
					if (sko='1') then
						if f_com= "00" then
							next_state <= s5;  -- для формата ПР  из s4 переходим в s5, если есть sko, запись младшей части результата в ОП
						else 
							next_state <= s0;	-- переходим в s0 для формата РР
						end if;
					else 	
						next_state <= s4; -- ждем завершения операции
					end if;
				when s5 =>
						next_state <= s6; -- Запись старшей части результата в ОП
				when s6 =>		
						next_state <= s0; -- из s6 всегда переходим в s0, это пустой такт, чтобы завершить запись в ОП и подать СК на адресный вход ОП,для выборки след ком
			end case;			
	end process NS;
---------------------------------------------------------------------------------------------------------
-- ниже приводится описание управляющих сигналов для БМК

incr_CK<='1' when (state=s0  or (state=s1 and f_com="00")) else -- разрешение на инкремент СК	всегда в s0  и в s1, если формат П-Р
			'0';
summ_CK<='1' when state=s1 and f_com="10" and priznak="10" else -- разрешение на приращение СК если выполняется условие перехода
			'0';
load_RK<='1' when (state=s0) else -- загрузка команды в RK всегда в s0 для любой операции
			'0';
load_RA<='1' when (state=s2) else -- загрузка ИА в RA в s2 для операции умножения
			'0';
incr_RA <='1' when (state=s4 and sko='1') else -- инкремент RA для записи старшей части результата в ОП, только для умножения
			'0';
sno <='1' when (state=s3) else -- когда извлекли операнды на шину А и В 
			'0';
wr_en_OP<='1' when ((state=s4 and sko='1' and f_com="00") or state=s5) else -- запись в ОП, если П-Р 
			'0';					
data_in_OP<= rr(2*n-1 downto n) when (state= s5) else
				 rr(n-1 downto 0);

address_OP <= CK	when (state=s0 or state=s1 or state=s6 or f_com="01") else -- если РР, то всегда CK
				  IA	when state=s2 else
				  RA; 
				  
IA<= data_out_OP+q_a; -- вычисляем исполнительный адрес первого операнда


wr_en_a_RP<='1' when state=s4 and sko='1' and f_com="01" else -- запись в РП, если формат Р-Р
				'0';

				
a<= data_out_OP when f_com="00" else --на шину А- первого операнда подаем первый операнд с выхода ОП, если формат память регистр
	 q_a;  -- 	либо с РП с выхода данных первого порта а, если формат регистр регистр 			  
b<= q_b; --на шину В - второго операнда подаем второй операнд, считанный через порт b РП	
 
-- сигнал f_com привязываем к полю сор, задаваемому в разрядах RK[7..6]
-- используем такое кодирование, как в восьмом проекте АУ: 00- сложение, 01-умножение
f_com<="00" when RK(7 downto 6)="01" else -- если умн, то ПР
		 "01" when RK(7 downto 6)="00" else -- если сложение, то РР
		 "10";		 -- если переход
		 
cop<=RK(6); -- этот разряд определяет операцию в арифметическом устройстве
---------------------------------------------------------------------------------------------------
wr_en_b_RP<='0'; --задаем в карте портов
address_a_RP<= RK (5 downto 3); -- поле R1  в команде
data_a_RP<= rr(7 downto 0); -- задаем в карте портов
address_b_RP<= RK (2 downto 0); -- поле R2  в команде, 
data_b_RP<= (others=>'0'); -- задаем все нули в карте портов
---------------------------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------
	--  отладочный выход для наблюдения текущего состояния
		s_out<="000" when state=s0 else
				  "001" when state=s1 else					
				  "010" when state=s2 else
				  "011" when state=s3 else
				  "100" when state=s4 else
				  "101" when state=s5 else
				  "110";
end arch;
